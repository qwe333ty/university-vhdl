library ieee;
use ieee.std_logic_1164.all;

-- Aliaksandr Rahavoi
entity test_entity is
end test_entity;

architecture test_architecture of test_entity is
    begin
end test_architecture;